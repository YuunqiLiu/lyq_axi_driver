AxiDriverSlave WriteMergeHandler need to support narrow transfer
Change all const to define value
Transaction length reduce
Interface X value process,Z/X和别的值做&&会被当做1