

module test();

    mailbox mbx;

    initial begin

    $display("$d",3/2);


    end



endmodule 