

class driver();


endclass