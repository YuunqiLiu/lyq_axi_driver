`define AXI_IF_AWID_WIDTH   32
`define AXI_IF_AWADDR_WIDTH 64
`define AXI_IF_AWLEN_WIDTH  4
`define AXI_IF_WID_WIDTH    32
`define AXI_IF_WDATA_WIDTH  1024
`define AXI_IF_WSTRB_WIDTH  128
`define AXI_IF_BID_WIDTH    32
`define AXI_IF_ARID_WIDTH   32
`define AXI_IF_ARADDR_WIDTH 64
`define AXI_IF_ARLEN_WIDTH  4
`define AXI_IF_RID_WIDTH    32
`define AXI_IF_RDATA_WIDTH  1024

`define AXI_IF_MASTER_NUM   16
`define AXI_IF_SLAVE_NUM    16
`define AXI_IF_MONITOR_NUM  16