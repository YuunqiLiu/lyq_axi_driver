
class AxiWChannelDataPack;

    bit [7:0]       data[4095:0];
    bit             strb[4095:0];
    bit [127:0]     user[255:0];

endclass